class spi_base_test extends uvm_test;
  `uvm_component_utils(spi_base_test)

  spi_env env;
  spi_seq seq;

  function new(string name, uvm_component parent);
    super.new(name, parent);
  endfunction

  function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    env = spi_env::type_id::create("env", this);
  endfunction

  task run_phase(uvm_phase phase);
    seq = spi_seq::type_id::create("seq");

    phase.raise_objection(this);
    `uvm_info("BASE_TEST", "Base test running", UVM_LOW)

    fork
      seq.start(env.agt.sqr);

    join

    phase.drop_objection(this);
  endtask
endclass