// Lets say that the environment class was already there, and generator is
// a new component that needs to be included in the ENV.
class env #( int LOOP, int ADDR_WIDTH, int DATA_WIDTH, bit [ADDR_WIDTH-1:0] ADDR_DIV );
  generator 	    #(.LOOP(LOOP), .ADDR_WIDTH(ADDR_WIDTH), .DATA_WIDTH(DATA_WIDTH))	        g0; 			// Generate transactions
  driver 			#(.ADDR_WIDTH(ADDR_WIDTH), .DATA_WIDTH(DATA_WIDTH))                         d0; 			// Driver to design
  monitor 		    #(.ADDR_WIDTH(ADDR_WIDTH), .DATA_WIDTH(DATA_WIDTH))                         m0_in; 			// Monitor driver to design
  monitor 		    #(.ADDR_WIDTH(ADDR_WIDTH), .DATA_WIDTH(DATA_WIDTH))                         m0_out; 	    // Monitor design to scoreboard
  scoreboard 		#(.ADDR_WIDTH(ADDR_WIDTH), .DATA_WIDTH(DATA_WIDTH), .ADDR_DIV(ADDR_DIV))    s0; 			// Scoreboard connected to monitor
  virtual switch_if #(.ADDR_WIDTH(ADDR_WIDTH), .DATA_WIDTH(DATA_WIDTH))                         m_switch_vif_in; 	// Virtual interface handle inputs
  virtual switch_if #(.ADDR_WIDTH(ADDR_WIDTH), .DATA_WIDTH(DATA_WIDTH))                         m_switch_vif_out; 	// Virtual interface handle outputs
  virtual clk_if 	                                                                            m_clk_vif; 		// TB clk

  event drv_done;
  mailbox drv_mbx, scb_mbx_in, scb_mbx_out;
  // mailbox scb_mbx; 		// Top level mailbox for SCB <-> MON

  function new();
    $display("T=%0t [Env] constructor", $time);
    d0 = new();
    m0_in = new();
    m0_out = new();
    s0 = new();
    // scb_mbx = new();
    g0 = new();
    drv_mbx = new();
    scb_mbx_in = new();
    scb_mbx_out = new();
  endfunction

  virtual task run();
    $display("T=%0t [Env] run task", $time);

    // Connect virtual interface handles
    d0.m_switch_vif = m_switch_vif_in;
    m0_in.m_switch_vif = m_switch_vif_in;
    m0_out.m_switch_vif = m_switch_vif_out;
    d0.m_clk_vif = m_clk_vif;
    m0_in.m_clk_vif = m_clk_vif;
    m0_out.m_clk_vif = m_clk_vif;

    // Connect mailboxes between each component
    d0.drv_mbx = drv_mbx;
    g0.drv_mbx = drv_mbx;

    // Mailboxes for input/output of scoreboard
    s0.scb_mbx_in = scb_mbx_in;
    m0_in.scb_mbx = scb_mbx_in;
    s0.scb_mbx_out = scb_mbx_out;
    m0_out.scb_mbx = scb_mbx_out;

    // Connect event handles
    d0.drv_done = drv_done;
    g0.drv_done = drv_done;

    // Start all components - a fork join_any is used because
    // the stimulus is generated by the generator and we want the
    // simulation to exit only when the generator has finished
    // creating all transactions. Until then all other components
    // have to run in the background.

    $display("T=%0t [Env] to start fork", $time);

    fork
    	s0.run();
		d0.run();
    	m0_in.run();
    	m0_out.run();
      	g0.run();
    join_any
  endtask
endclass
