class fa_test extends uvm_test;
  `uvm_component_utils(fa_test)

  fa_env env;

  function new(string name, uvm_component parent);
    super.new(name, parent);
  endfunction

  function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    env = fa_env::type_id::create("env", this);
  endfunction

endclass
