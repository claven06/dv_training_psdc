// This is a one-line comment

/* This is a multiple line comment.
Since this line is within the block comment symbols, it is a comment.
*/

/* Another multiple line comment
// A nested one-line comment inside a block comment is fine.
But a block comment cannot be nested in another block comment.
*/
