package ptop_uvm_pkg;

  // Re-export all sub-packages
  import ptop_child_pkg::*;
  import ptop_parent_pkg::*; 
  import ptop_test_pkg::*;

endpackage
